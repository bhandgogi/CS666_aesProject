module SubTable(state, stateOut);
	input [7:0] state; // Original byte
	output reg [7:0] stateOut; // Corresponding sub_byte
    
	always @(state) begin
		case (state)
			8'h00: stateOut=8'h63;
			8'h01: stateOut=8'h7c;
			8'h02: stateOut=8'h77;
			8'h03: stateOut=8'h7b;
			8'h04: stateOut=8'hf2;
			8'h05: stateOut=8'h6b;
			8'h06: stateOut=8'h6f;
			8'h07: stateOut=8'hc5;
			8'h08: stateOut=8'h30;
			8'h09: stateOut=8'h01;
			8'h0a: stateOut=8'h67;
			8'h0b: stateOut=8'h2b;
			8'h0c: stateOut=8'hfe;
			8'h0d: stateOut=8'hd7;
			8'h0e: stateOut=8'hab;
			8'h0f: stateOut=8'h76;
			8'h10: stateOut=8'hca;
			8'h11: stateOut=8'h82;
			8'h12: stateOut=8'hc9;
			8'h13: stateOut=8'h7d;
			8'h14: stateOut=8'hfa;
			8'h15: stateOut=8'h59;
			8'h16: stateOut=8'h47;
			8'h17: stateOut=8'hf0;
			8'h18: stateOut=8'had;
			8'h19: stateOut=8'hd4;
			8'h1a: stateOut=8'ha2;
			8'h1b: stateOut=8'haf;
			8'h1c: stateOut=8'h9c;
			8'h1d: stateOut=8'ha4;
			8'h1e: stateOut=8'h72;
			8'h1f: stateOut=8'hc0;
			8'h20: stateOut=8'hb7;
			8'h21: stateOut=8'hfd;
			8'h22: stateOut=8'h93;
			8'h23: stateOut=8'h26;
			8'h24: stateOut=8'h36;
			8'h25: stateOut=8'h3f;
			8'h26: stateOut=8'hf7;
			8'h27: stateOut=8'hcc;
			8'h28: stateOut=8'h34;
			8'h29: stateOut=8'ha5;
			8'h2a: stateOut=8'he5;
			8'h2b: stateOut=8'hf1;
			8'h2c: stateOut=8'h71;
			8'h2d: stateOut=8'hd8;
			8'h2e: stateOut=8'h31;
			8'h2f: stateOut=8'h15;
			8'h30: stateOut=8'h04;
			8'h31: stateOut=8'hc7;
			8'h32: stateOut=8'h23;
			8'h33: stateOut=8'hc3;
			8'h34: stateOut=8'h18;
			8'h35: stateOut=8'h96;
			8'h36: stateOut=8'h05;
			8'h37: stateOut=8'h9a;
			8'h38: stateOut=8'h07;
			8'h39: stateOut=8'h12;
			8'h3a: stateOut=8'h80;
			8'h3b: stateOut=8'he2;
			8'h3c: stateOut=8'heb;
			8'h3d: stateOut=8'h27;
			8'h3e: stateOut=8'hb2;
			8'h3f: stateOut=8'h75;
			8'h40: stateOut=8'h09;
			8'h41: stateOut=8'h83;
			8'h42: stateOut=8'h2c;
			8'h43: stateOut=8'h1a;
			8'h44: stateOut=8'h1b;
			8'h45: stateOut=8'h6e;
			8'h46: stateOut=8'h5a;
			8'h47: stateOut=8'ha0;
			8'h48: stateOut=8'h52;
			8'h49: stateOut=8'h3b;
			8'h4a: stateOut=8'hd6;
			8'h4b: stateOut=8'hb3;
			8'h4c: stateOut=8'h29;
			8'h4d: stateOut=8'he3;
			8'h4e: stateOut=8'h2f;
			8'h4f: stateOut=8'h84;
			8'h50: stateOut=8'h53;
			8'h51: stateOut=8'hd1;
			8'h52: stateOut=8'h00;
			8'h53: stateOut=8'hed;
			8'h54: stateOut=8'h20;
			8'h55: stateOut=8'hfc;
			8'h56: stateOut=8'hb1;
			8'h57: stateOut=8'h5b;
			8'h58: stateOut=8'h6a;
			8'h59: stateOut=8'hcb;
			8'h5a: stateOut=8'hbe;
			8'h5b: stateOut=8'h39;
			8'h5c: stateOut=8'h4a;
			8'h5d: stateOut=8'h4c;
			8'h5e: stateOut=8'h58;
			8'h5f: stateOut=8'hcf;
			8'h60: stateOut=8'hd0;
			8'h61: stateOut=8'hef;
			8'h62: stateOut=8'haa;
			8'h63: stateOut=8'hfb;
			8'h64: stateOut=8'h43;
			8'h65: stateOut=8'h4d;
			8'h66: stateOut=8'h33;
			8'h67: stateOut=8'h85;
			8'h68: stateOut=8'h45;
			8'h69: stateOut=8'hf9;
			8'h6a: stateOut=8'h02;
			8'h6b: stateOut=8'h7f;
			8'h6c: stateOut=8'h50;
			8'h6d: stateOut=8'h3c;
			8'h6e: stateOut=8'h9f;
			8'h6f: stateOut=8'ha8;
			8'h70: stateOut=8'h51;
			8'h71: stateOut=8'ha3;
			8'h72: stateOut=8'h40;
			8'h73: stateOut=8'h8f;
			8'h74: stateOut=8'h92;
			8'h75: stateOut=8'h9d;
			8'h76: stateOut=8'h38;
			8'h77: stateOut=8'hf5;
			8'h78: stateOut=8'hbc;
			8'h79: stateOut=8'hb6;
			8'h7a: stateOut=8'hda;
			8'h7b: stateOut=8'h21;
			8'h7c: stateOut=8'h10;
			8'h7d: stateOut=8'hff;
			8'h7e: stateOut=8'hf3;
			8'h7f: stateOut=8'hd2;
			8'h80: stateOut=8'hcd;
			8'h81: stateOut=8'h0c;
			8'h82: stateOut=8'h13;
			8'h83: stateOut=8'hec;
			8'h84: stateOut=8'h5f;
			8'h85: stateOut=8'h97;
			8'h86: stateOut=8'h44;
			8'h87: stateOut=8'h17;
			8'h88: stateOut=8'hc4;
			8'h89: stateOut=8'ha7;
			8'h8a: stateOut=8'h7e;
			8'h8b: stateOut=8'h3d;
			8'h8c: stateOut=8'h64;
			8'h8d: stateOut=8'h5d;
			8'h8e: stateOut=8'h19;
			8'h8f: stateOut=8'h73;
			8'h90: stateOut=8'h60;
			8'h91: stateOut=8'h81;
			8'h92: stateOut=8'h4f;
			8'h93: stateOut=8'hdc;
			8'h94: stateOut=8'h22;
			8'h95: stateOut=8'h2a;
			8'h96: stateOut=8'h90;
			8'h97: stateOut=8'h88;
			8'h98: stateOut=8'h46;
			8'h99: stateOut=8'hee;
			8'h9a: stateOut=8'hb8;
			8'h9b: stateOut=8'h14;
			8'h9c: stateOut=8'hde;
			8'h9d: stateOut=8'h5e;
			8'h9e: stateOut=8'h0b;
			8'h9f: stateOut=8'hdb;
			8'ha0: stateOut=8'he0;
			8'ha1: stateOut=8'h32;
			8'ha2: stateOut=8'h3a;
			8'ha3: stateOut=8'h0a;
			8'ha4: stateOut=8'h49;
			8'ha5: stateOut=8'h06;
			8'ha6: stateOut=8'h24;
			8'ha7: stateOut=8'h5c;
			8'ha8: stateOut=8'hc2;
			8'ha9: stateOut=8'hd3;
			8'haa: stateOut=8'hac;
			8'hab: stateOut=8'h62;
			8'hac: stateOut=8'h91;
			8'had: stateOut=8'h95;
			8'hae: stateOut=8'he4;
			8'haf: stateOut=8'h79;
			8'hb0: stateOut=8'he7;
			8'hb1: stateOut=8'hc8;
			8'hb2: stateOut=8'h37;
			8'hb3: stateOut=8'h6d;
			8'hb4: stateOut=8'h8d;
			8'hb5: stateOut=8'hd5;
			8'hb6: stateOut=8'h4e;
			8'hb7: stateOut=8'ha9;
			8'hb8: stateOut=8'h6c;
			8'hb9: stateOut=8'h56;
			8'hba: stateOut=8'hf4;
			8'hbb: stateOut=8'hea;
			8'hbc: stateOut=8'h65;
			8'hbd: stateOut=8'h7a;
			8'hbe: stateOut=8'hae;
			8'hbf: stateOut=8'h08;
			8'hc0: stateOut=8'hba;
			8'hc1: stateOut=8'h78;
			8'hc2: stateOut=8'h25;
			8'hc3: stateOut=8'h2e;
			8'hc4: stateOut=8'h1c;
			8'hc5: stateOut=8'ha6;
			8'hc6: stateOut=8'hb4;
			8'hc7: stateOut=8'hc6;
			8'hc8: stateOut=8'he8;
			8'hc9: stateOut=8'hdd;
			8'hca: stateOut=8'h74;
			8'hcb: stateOut=8'h1f;
			8'hcc: stateOut=8'h4b;
			8'hcd: stateOut=8'hbd;
			8'hce: stateOut=8'h8b;
			8'hcf: stateOut=8'h8a;
			8'hd0: stateOut=8'h70;
			8'hd1: stateOut=8'h3e;
			8'hd2: stateOut=8'hb5;
			8'hd3: stateOut=8'h66;
			8'hd4: stateOut=8'h48;
			8'hd5: stateOut=8'h03;
			8'hd6: stateOut=8'hf6;
			8'hd7: stateOut=8'h0e;
			8'hd8: stateOut=8'h61;
			8'hd9: stateOut=8'h35;
			8'hda: stateOut=8'h57;
			8'hdb: stateOut=8'hb9;
			8'hdc: stateOut=8'h86;
			8'hdd: stateOut=8'hc1;
			8'hde: stateOut=8'h1d;
			8'hdf: stateOut=8'h9e;
			8'he0: stateOut=8'he1;
			8'he1: stateOut=8'hf8;
			8'he2: stateOut=8'h98;
			8'he3: stateOut=8'h11;
			8'he4: stateOut=8'h69;
			8'he5: stateOut=8'hd9;
			8'he6: stateOut=8'h8e;
			8'he7: stateOut=8'h94;
			8'he8: stateOut=8'h9b;
			8'he9: stateOut=8'h1e;
			8'hea: stateOut=8'h87;
			8'heb: stateOut=8'he9;
			8'hec: stateOut=8'hce;
			8'hed: stateOut=8'h55;
			8'hee: stateOut=8'h28;
			8'hef: stateOut=8'hdf;
			8'hf0: stateOut=8'h8c;
			8'hf1: stateOut=8'ha1;
			8'hf2: stateOut=8'h89;
			8'hf3: stateOut=8'h0d;
			8'hf4: stateOut=8'hbf;
			8'hf5: stateOut=8'he6;
			8'hf6: stateOut=8'h42;
			8'hf7: stateOut=8'h68;
			8'hf8: stateOut=8'h41;
			8'hf9: stateOut=8'h99;
			8'hfa: stateOut=8'h2d;
			8'hfb: stateOut=8'h0f;
			8'hfc: stateOut=8'hb0;
			8'hfd: stateOut=8'h54;
			8'hfe: stateOut=8'hbb;
			8'hff: stateOut=8'h16;
		endcase
	end
endmodule